module ex19_top();

endmodule
